`timescale 1ns/1ns
module UnidadDeControl (input [5:0] InstruccionControl, output RegDst, output Branch, output MemToReg, output [3:0] ALUOp, output ALUSrc, output RegWrite);

endmodule
