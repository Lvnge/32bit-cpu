`timescale 1ns/1ns
module Alucontrol (input [5:0] inst, input [3:0] ALUOp, output [2:0] instalu);

endmodule
